`timescale 1 ps / 1 ps

module IOBUFDS_DCIEN_model #(
  parameter IBUF_LOW_PWR = "TRUE",
  parameter SLEW = "SLOW",
  parameter USE_IBUFDISABLE = "TRUE"
)(
  output O,
  inout IO,
  inout IOB,
  input DCITERMDISABLE,
  input I,
  input IBUFDISABLE,
  input T
);
 // black box
endmodule
