`timescale  1 ps / 1 ps

module IOBUF_DCIEN_model #(
  parameter IBUF_LOW_PWR = "TRUE",
  parameter SLEW = "SLOW",
  parameter USE_IBUFDISABLE = "TRUE"
)(
  output O,
  inout IO,
  input I,
  input T,
  input DCITERMDISABLE,
  input IBUFDISABLE
);
// black box

endmodule

